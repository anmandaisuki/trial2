module xor ();

assign a = 1'b0;