module xor ();